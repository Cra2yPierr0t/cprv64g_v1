module cprv_rom_1p #(
    parameter ADDR_WIDTH    = 7,
    parameter DATA_WIDTH    = 64
)(
    input   logic                  clk,
    input   logic                  w_en,
    input   logic [ADDR_WIDTH-1:0] addr,
    input   logic [DATA_WIDTH-1:0] wdata,
    output  logic [DATA_WIDTH-1:0] rdata
);

    logic [DATA_WIDTH-1:0] mem [2**ADDR_WIDTH-1:0];

    always_ff @(posedge clk) begin
        if(w_en) begin
            mem[addr >> 2] <= wdata;
            rdata <= wdata;
        end else begin
            rdata <= mem[addr >> 2];
        end
    end

    integer i;
    initial begin
        mem[0] = 32'b000000000001_00001_000_00001_0010011;
        mem[1] = 32'b000000000001_00001_000_00001_0010011;
        mem[2] = 32'b000000000001_00001_000_00001_0010011;
        mem[3] = 32'b000000000001_00001_000_00001_0010011;
        mem[4] = 32'b000000000001_00001_000_00001_0010011;
        mem[5] = 32'b000000000001_00001_000_00001_0010011;
        mem[6] = 32'b000000000001_00001_000_00001_0010011;
        mem[7] = 32'b000000000001_00001_000_00001_0010011;
        mem[8] = 32'b000000000001_00001_000_00001_0010011;
        mem[9] = 32'b000000000001_00001_000_00001_0010011;
        mem[10] = 32'b000000000001_00001_000_00001_0010011;
        mem[11] = 32'b000000000001_00001_000_00001_0010011;

        mem[12] = 32'b0000000_00001_00000_010_00000_0100011;
        mem[13] = 32'b0000000_00001_00000_010_00000_0100011;
        mem[14] = 32'b0000000_00001_00000_010_00000_0100011;
        mem[15] = 32'b0000000_00001_00000_010_00000_0100011;
        mem[16] = 32'b0000000_00001_00000_010_00000_0100011;
        mem[17] = 32'b000000000001_00000_010_00010_0000011;
    end

endmodule
