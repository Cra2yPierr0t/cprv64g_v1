module cprv_sim (
    input logic clk
);

    cprv_top top (
        .clk    (clk    )
    );
endmodule
